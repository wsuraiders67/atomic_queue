-- _____________________________________________________________________________
--|
--|      sssssssss     nnnn nnnnnnn      cccccccccc
--|     sssssssssss    nnnnn    nnnn    cccccccccccc
--|     ssss   ssss    nnnn     nnnn    cccc    cccc    Sierra
--|     ssss           nnnn     nnnn    cccc    cccc    Nevada
--|      sssssssss     nnnn     nnnn    cccc            Corporation
--|            ssss    nnnn     nnnn    cccc    cccc
--|     ssss   ssss    nnnn     nnnn    cccc    cccc
--|     sssssssssss    nnnn     nnnn    cccccccccccc
--|      sssssssss     nnnn     nnnn     cccccccccc     Copyright 2015
--|_____________________________________________________________________________
--|
--|      //  //======  Sensor Systems and Technologies
--|     ||  ||   ||    2611 Commons Blvd
--|      \\  \\  ||    Beavercreek, OH 45431
--|       ||  || ||
--|      //  //  ||    937-431-2800
--|_____________________________________________________________________________
--|
--|       File              : axi_pkg
--|       Original Project  : GS Maven
--|       Original Author   : Craig McGillivary
--|       Original Date     : 8/22/2019
--|_____________________________________________________________________________
--|
--|     Description : Definitions (records, etc.) for AXI-4 Lite interfaces
--|     Information was gathered from "AMBA AXI and ACE Protocol Specification"
--|     copyright 2003 ARM
--|
--|   The AXI specification defines several types of busses, of 2 different directions.
--| There is a "command" record that's generated by the AXI Master to request reads or
--| writes of the AXI Slave devices on the bus. The Slave devices then generate a
--| "response" record that contains the results of the read or write.
--|   The AXI Lite bus is the simplest of all, and transfers a single value
--| during each transaction. This package contains the definitions of the AXI Lite
--| records. (Again that's a command record from the Master, and a response record
--| from the Slave.) The at its simplist AXIL uses 32 address bits and 32 data bits
--| but it can use up to 64 address and 64 data.
--|   The AXI Stream allows multiple and individual bytes to be transferred "on demand"
--| and without the overhead associated with providing addresses.  All of the response
--| records for AXI streams are really the same type with different aliases since the
--| record only includes a tready signal.
--|   The full-up AXI bus (aka AXI Memory Mapped) is the most complicated and can
--| transfer bursts of variable sized data during each transaction. Plus it can use
--| 32-bit or 64-bit addresses.
--|   Conversion between axi packages of different data widths is not recommended.
--| However converting axi command records from one address width to another can be
--| done by using overloaded axi_addr_resize functions. Converting axi response
--| records for different address widths is easier because the records have no
--| address members. We actually use aliases so rt_axil32x64_rsp and axil_rsp are
--| really the same object and no conversion function is needed for response records
--| as long as the data widths are the same.
--|   It is recommended that for full axi records you use the 64 bit address version
--| and then leave the upper bits unconnected. A similar style is recommended for ID
--| bits since the number of ID bits carried through different parts of the
--| interconnect grows and it is better not to have lots of different AXI types.
--|
--|
--|   The AXI records defined in the entity are:
--|     -- AXI Lites
--|       rt_axil_cmd       -- AXI Lite "command" record from the Master to the Slave, 32 bit data path, 32 bit address
--|       rt_axil_rsp       -- AXI Lite "response" record from the Slave to the Master 32 bit data path, 32 bit address
--|       rt_axil32x16_cmd  -- AXI Lite "command" record from the Master to the Slave, 32 bit data path, 16 bit address
--|       rt_axil32x16_rsp  -- AXI Lite "response" record from the Slave to the Master 32 bit data path, 16 bit address
--|       rt_axil32x64_cmd  -- same as above, but with a 32 bit data path, 64 bit address
--|       rt_axil32x64_rsp
--|       rt_axil64x32_cmd  -- same as above, but with a 64 bit data path, 32 bit address
--|       rt_axil64x32_rsp
--|       rt_axil64x40_cmd  -- same as above, but with a 64 bit data path, 40 bit address
--|       rt_axil64x40_rsp
--|       rt_axil64x64_cmd  -- same as above, but with a 64 bit data path, 64 bit address
--|       rt_axil64x64_rsp
--|
--|     -- AXI Streams
--|       rt_axis16_cmd     -- AXI Stream command record from the Master, 32 bit wide data path
--|       rt_axis16_rsp     -- AXI Stream response record from the Slave
--|       rt_axis32_cmd     -- AXI Stream command record from the Master, 32 bit wide data path
--|       rt_axis32_rsp     -- AXI Stream response record from the Slave
--|       rt_axis64_cmd     -- same as above, but with a 64 bit wide data path
--|       rt_axis64_rsp
--|       rt_axis128_cmd    -- same as above, but with a 128 bit wide data path
--|       rt_axis128_rsp
--|       rt_axis256_cmd    -- same as above, but with a 256 bit wide data path
--|       rt_axis256_rsp
--|       rt_axis512_cmd    -- same as above, but with a 512 bit wide data path
--|       rt_axis512_rsp
--|       rt_axis1024_cmd    -- same as above, but with a 1024 bit wide data path
--|       rt_axis1024_rsp
--|
--|     -- Full AXI4 (aka AXI Memory Mapped)
--|       -- legacy 32 bit address records
--|       rt_axi32x32_cmd   -- AXI "command" record from the Master to the Slave, 32 bit data path, 32 bit address
--|       rt_axi32x32_rsp   -- AXI "response" record from the Slave to the Master 32 bit data path  32 bit address
--|       rt_axi64x32_cmd   -- same as above, but with a  64 bit data path, 32 bit address
--|       rt_axi64x32_rsp
--|       rt_axi64x32x16_cmd -- same as above, but with 16-bit ID
--|       rt_axi64x32x16_rsp
--|       rt_axi512x32_cmd  -- same as above, but with a  512 bit data path, 32 bit address
--|       rt_axi512x32_rsp
--|       rt_axi_mpsoc64_cmd-- same as above, but with a  64 bit data path, 40 bit address
--|       rt_axi_mpsoc64_rsp
--|       rt_axi_mpsoc32_cmd-- same as above, but with a  32 bit data path, 40 bit address
--|       rt_axi_mpsoc32_rsp
--|       rt_axi32_cmd      -- same as above, but with a   32 bit data path, 64 bit address
--|       rt_axi32_rsp
--|       rt_axi64_cmd      -- same as above, but with a   64 bit data path, 64 bit address
--|       rt_axi64_rsp
--|       rt_axi128_cmd     -- same as above, but with a  128 bit data path, 64 bit address
--|       rt_axi128_rsp
--|       rt_axi256_cmd     -- same as above, but with a  256 bit data path, 64 bit address
--|       rt_axi256_rsp
--|       rt_axi512_cmd     -- same as above, but with a  512 bit data path, 64 bit address
--|       rt_axi512_rsp
--|       rt_axi1024_cmd    -- same as above, but with a 1024 bit data path, 64 bit address
--|       rt_axi1024_rsp
--|
--|     -- Overloaded functions to change AXI command records to/from 64 bit addressing
--|       axi_addr_resize   -- go from 64 bit addressing to 32 bit addressing or the opposite
--|
--|   NOTE: The naming convention is:
--|     "axil" is an AXI Lite 32 data bits and 32 address bits,
--|     "axisXX" is an AXI Stream with an XX bit wide data path
--|     "axiXX" is a full-up AXI Memory Map with an XX bit wide data path abd 64 bit address bits
--      "axiDDxAA" is a full-up AXI Memory Map with an DD bit wide data path abd AA bit address bits
--|
--+-----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package axi_pkg is

  --************************************************************************
  --
  --    These enumerated types declare the possible burst sizes, as specified
  -- in either awsize or arsize.
  --
  --************************************************************************
  constant E_SIZE_001BYTES    : std_logic_vector(2 downto 0) := "000";
  constant E_SIZE_002BYTES    : std_logic_vector(2 downto 0) := "001";
  constant E_SIZE_004BYTES    : std_logic_vector(2 downto 0) := "010";
  constant E_SIZE_008BYTES    : std_logic_vector(2 downto 0) := "011";
  constant E_SIZE_016BYTES    : std_logic_vector(2 downto 0) := "100";
  constant E_SIZE_032BYTES    : std_logic_vector(2 downto 0) := "101";
  constant E_SIZE_064BYTES    : std_logic_vector(2 downto 0) := "110";
  constant E_SIZE_128BYTES    : std_logic_vector(2 downto 0) := "111";

  --************************************************************************
  --
  --    Here are the enumerated types of bursts, as specified by either awburst
  -- or arburst fields. The burst type and the size information, determine how
  -- the address for each transfer within the burst is calculated.
  --
  --************************************************************************
  constant E_BURST_FIXED      : std_logic_vector(1 downto 0) := "00";       -- Multiple reads or writes to the same address
  constant E_BURST_INCR       : std_logic_vector(1 downto 0) := "01";       -- Address increments by 2^awsize or 2^arsize
  constant E_BURST_WRAP       : std_logic_vector(1 downto 0) := "10";       -- Similar to INCR but will wrap at an address boundary

  --************************************************************************
  --
  --    The Lock type is specified for either awlock or arlock. It provides
  -- additional info about the atomic characteristics of the transfer.
  --
  --************************************************************************
  constant E_LOCK_NORM        : std_logic_vector(0 downto 0) := "0";        -- Normal access
  constant E_LOCK_EXLUSIVE    : std_logic_vector(0 downto 0) := "1";        -- Exclusive Access

  --************************************************************************
  --
  --    These enumerated types are the possible responses as specified by either
  -- rresp or bresp.
  --
  --************************************************************************
  constant E_RESP_OKAY        : std_logic_vector(1 downto 0) := "00";       -- Normal access success, or can indicate exclusive access failed
  constant E_RESP_EXOKAY      : std_logic_vector(1 downto 0) := "01";       -- Exclusive access has been successful
  constant E_RESP_SLVERR      : std_logic_vector(1 downto 0) := "10";       -- Slave error, the slave wishes to return an error master
  constant E_RESP_DECERR      : std_logic_vector(1 downto 0) := "11";       -- Decode error (by an interconnect component), no slave at addr

  --************************************************************************
  --
  --   This enumeration type is the the Xilinx recommended values for AWCACHE
  -- and ARCACHE. These are the values used by all Xilinx IP and recommended
  -- by the AXI Reference Guide UG761.
  --
  --************************************************************************
  constant E_NORM_NCACH_MOD_BUF : std_logic_vector(3 downto 0) := "0011";   --Normal, Non-cacheable, Modifiable and Bufferable

  --************************************************************************
  --
  --   This enumeration type is the the Xilinx recommended values for AWPROT
  -- and ARPROT. These are the values used by all Xilinx IP and recommended
  -- by the AXI Reference Guide UG761.
  --
  --************************************************************************
  constant E_NORM_SEC_DATA    : std_logic_vector(2 downto 0) := "000";      --Normal, Secure and Data

  --************************************************************************
  --
  --    Record for AXI4 Lite commands. This record contains all the signals
  -- sourced by the Master (the master initiates all transactions on the bus).
  -- These signals are grouped into 5 unique channels as specified by the AXI4
  -- protocol.
  --    The constant is used to zero-out unconnected rt_axil_cmd signals. If left
  -- unconnected, an axi interface could lock up because it is waiting for a
  -- "valid" signal.
  --
  --************************************************************************
  type rt_axil_cmd is
  record
    -- Write Address Channel Signals
    awaddr    : std_logic_vector(31 downto 0);    -- Write address gives the address of the single transfer
    awcache   : std_logic_vector( 3 downto 0);    -- Memory type indicates how transactions progress through a system
    awprot    : std_logic_vector( 2 downto 0);    -- Protection type indicates the privilege and security level
    awvalid   : std_logic;                        -- Write address valid, the channel is signaling address and control information
    -- Write Data Channel Signals
    wdata     : std_logic_vector(31 downto 0);    -- Xilinx documentation states the AXI4-Lite does not support 64 bit data 2012/01/18
    wstrb     : std_logic_vector( 3 downto 0);    -- Write strobes indicate which byte lanes (in wdata) hold valid data
    wvalid    : std_logic;                        -- Write valid indicates that write data and strobes are available
    -- Write Response Channel
    bready    : std_logic;                        -- Response ready indicates that the master can accept a write response
    -- Read Address Channel
    araddr    : std_logic_vector(31 downto 0);    -- Read address gives the address of the single transfer
    arcache   : std_logic_vector( 3 downto 0);    -- Memory type indicates how transactions progress through a system
    arprot    : std_logic_vector( 2 downto 0);    -- Protection type, privilege and security level of the transaction
    arvalid   : std_logic;                        -- Read address valid, the channel is signaling address and control information
    -- Read Data Channel
    rready    : std_logic;                        -- Read ready indicates the master can accept a read response
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL_CMD_RST     : rt_axil_cmd := (
    awaddr    => (others => '0'),
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wvalid    => '0',
    bready    => '0',
    araddr    => (others => '0'),
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arvalid   => '0',
    rready    => '0'
    );

  type at_axil_cmd is array (natural range <>) of rt_axil_cmd;

  --************************************************************************
  --
  --    Record for AXI4 Lite responses. This record contains all the signals
  -- sourced by the Slave (the slave responds to transactions on the bus).
  -- These signals are grouped into 5 unique channels as specified by the AXI4
  -- protocol.
  --    The constant is used to zero-out unconnected rt_axil_rsp signals. If left
  -- unconnected, an axi interface could lock up because it is waiting for a
  -- "valid" signal.
  --
  --************************************************************************
  type rt_axil_rsp is
  record
    -- Write Address Channel Signals
    awready   : std_logic;                        -- Write address ready, the slave is ready to accept an address and control signals
    -- Write Data Channel Signals
    wready    : std_logic;                        -- Write ready indicates that the slave can accept the write data
    -- Write Response Channel
    bresp     : std_logic_vector( 1 downto 0);    -- Xilinx documentation states the AXI4-Lite does not support EXOKAY response 2012/01/18
    bvalid    : std_logic;                        -- Write response valid indicates that the channel is signaling a valid write response
    -- Read Address Channel
    arready   : std_logic;                        -- Read address ready, the slave is ready to accept an address and control signals
    -- Read Data Channel
    rdata     : std_logic_vector(31 downto 0);    -- Xilinx documentation states the AXI4-Lite does not support 64 bit data 2012/01/18
    rresp     : std_logic_vector( 1 downto 0);    -- Xilinx documentation states the AXI4-Lite does not support EXOKAY response 2012/01/18
    rvalid    : std_logic;                        -- Read valid indicates the channel is signaling the requested read data
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL_RSP_RST     : rt_axil_rsp := (
    awready   => '0',
    wready    => '0',
    bresp     => E_RESP_OKAY,
    bvalid    => '0',
    arready   => '0',
    rdata     => (others => '0'),
    rresp     => E_RESP_OKAY,
    rvalid    => '0'
    );

  type at_axil_rsp is array (natural range <>) of rt_axil_rsp;

  --************************************************************************
  --
  --    AXI Lite command for 32- bit data path and 16 bit addresses.
  --
  --************************************************************************
  type rt_axil32x16_cmd is
  record
    -- Write Address Channel Signals
    awaddr    : std_logic_vector(15 downto 0);    -- Write address gives the address of the single transfer
    awcache   : std_logic_vector( 3 downto 0);    -- Memory type indicates how transactions progress through a system
    awprot    : std_logic_vector( 2 downto 0);    -- Protection type indicates the privilege and security level
    awvalid   : std_logic;                        -- Write address valid, the channel is signaling address and control information
    -- Write Data Channel Signals
    wdata     : std_logic_vector(31 downto 0);    -- Xilinx documentation states the AXI4-Lite does not support 64 bit data 2012/01/18
    wstrb     : std_logic_vector( 3 downto 0);    -- Write strobes indicate which byte lanes (in wdata) hold valid data
    wvalid    : std_logic;                        -- Write valid indicates that write data and strobes are available
    -- Write Response Channel
    bready    : std_logic;                        -- Response ready indicates that the master can accept a write response
    -- Read Address Channel
    araddr    : std_logic_vector(15 downto 0);    -- Read address gives the address of the single transfer
    arcache   : std_logic_vector( 3 downto 0);    -- Memory type indicates how transactions progress through a system
    arprot    : std_logic_vector( 2 downto 0);    -- Protection type, privilege and security level of the transaction
    arvalid   : std_logic;                        -- Read address valid, the channel is signaling address and control information
    -- Read Data Channel
    rready    : std_logic;                        -- Read ready indicates the master can accept a read response
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL32X16_CMD_RST     : rt_axil32x16_cmd := (
    awaddr    => (others => '0'),
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wvalid    => '0',
    bready    => '0',
    araddr    => (others => '0'),
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arvalid   => '0',
    rready    => '0'
    );

  type at_axil32x16_cmd is array (natural range <>) of rt_axil32x16_cmd;

  --************************************************************************
  --
  -- Even though there is no address bits in the response packets we can hide that
  -- detail from the user to make things clearer. We will use alias so that no
  -- conversion is needed between rt_axil_rsp and rt_axil32x64_rsp
  --
  --************************************************************************
  type rt_axil32x16_rsp is
  record
    -- Write Address Channel Signals
    awready   : std_logic;                        -- Write address ready, the slave is ready to accept an address and control signals
    -- Write Data Channel Signals
    wready    : std_logic;                        -- Write ready indicates that the slave can accept the write data
    -- Write Response Channel
    bresp     : std_logic_vector( 1 downto 0);    -- Xilinx documentation states the AXI4-Lite does not support EXOKAY response 2012/01/18
    bvalid    : std_logic;                        -- Write response valid indicates that the channel is signaling a valid write response
    -- Read Address Channel
    arready   : std_logic;                        -- Read address ready, the slave is ready to accept an address and control signals
    -- Read Data Channel
    rdata     : std_logic_vector(31 downto 0);    -- Xilinx documentation states the AXI4-Lite does not support 64 bit data 2012/01/18
    rresp     : std_logic_vector( 1 downto 0);    -- Xilinx documentation states the AXI4-Lite does not support EXOKAY response 2012/01/18
    rvalid    : std_logic;                        -- Read valid indicates the channel is signaling the requested read data
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL32X16_RSP_RST     : rt_axil32x16_rsp := (
    awready   => '0',
    wready    => '0',
    bresp     => E_RESP_OKAY,
    bvalid    => '0',
    arready   => '0',
    rdata     => (others => '0'),
    rresp     => E_RESP_OKAY,
    rvalid    => '0'
    );

  type at_axil32x16_rsp is array (natural range <>) of rt_axil32x16_rsp;

  --************************************************************************
  --
  --    AXI Lite command for 32- bit data path and  64 bit addresses.
  --
  --************************************************************************
  type rt_axil32x64_cmd is
  record
    -- Write Address Channel Signals
    awaddr    : std_logic_vector(63 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(31 downto 0);
    wstrb     : std_logic_vector( 3 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    araddr    : std_logic_vector(63 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL32x64_CMD_RST     : rt_axil32x64_cmd := (
    awaddr    => (others => '0'),
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wvalid    => '0',
    bready    => '0',
    araddr    => (others => '0'),
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arvalid   => '0',
    rready    => '0'
    );

  type at_axil32x64_cmd is array (natural range <>) of rt_axil32x64_cmd;

  --************************************************************************
  --
  -- Even though there is no address bits in the response packets we can hide that
  -- detail from the user to make things clearer. We will use alias so that no
  -- conversion is needed between rt_axil_rsp and rt_axil32x64_rsp
  --
  --************************************************************************
  alias rt_axil32x64_rsp    is rt_axil_rsp;
  alias K_AXIL32x64_RSP_RST is K_AXIL_RSP_RST;
  alias at_axil32x64_rsp    is at_axil_rsp;

  --************************************************************************
  --
  --    AXI Lite command for 64- bit data path and  32 bit addresses.
  --
  --************************************************************************
  type rt_axil64x32_cmd is
  record
    -- Write Address Channel Signals
    awaddr    : std_logic_vector(31 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(63 downto 0);
    wstrb     : std_logic_vector( 7 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    araddr    : std_logic_vector(31 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL64x32_CMD_RST     : rt_axil64x32_cmd := (
    awaddr    => (others => '0'),
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wvalid    => '0',
    bready    => '0',
    araddr    => (others => '0'),
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arvalid   => '0',
    rready    => '0'
    );

  type at_axil64x32_cmd is array (natural range <>) of rt_axil64x32_cmd;

  --************************************************************************
  --
  --    AXI Lite respone for 64- bit data path and  32 bit addresses.
  --
  --************************************************************************
  type rt_axil64x32_rsp is
  record
    -- Write Address Channel Signals
    awready   : std_logic;
    -- Write Data Channel Signals
    wready    : std_logic;
    -- Write Response Channel
    bresp     : std_logic_vector( 1 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rdata     : std_logic_vector(63 downto 0);
    rresp     : std_logic_vector( 1 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL64x32_RSP_RST     : rt_axil64x32_rsp := (
    awready   => '0',
    wready    => '0',
    bresp     => E_RESP_OKAY,
    bvalid    => '0',
    arready   => '0',
    rdata     => (others => '0'),
    rresp     => E_RESP_OKAY,
    rvalid    => '0'
    );

  type at_axil64x32_rsp is array (natural range <>) of rt_axil64x32_rsp;

  --************************************************************************
  --
  --    AXI Lite command for 64-bit data path and 40-bit addresses.
  --
  --************************************************************************
  type rt_axil64x40_cmd is
  record
    -- Write Address Channel Signals
    awaddr    : std_logic_vector(39 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(63 downto 0);
    wstrb     : std_logic_vector( 7 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    araddr    : std_logic_vector(39 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL64x40_CMD_RST     : rt_axil64x40_cmd := (
    awaddr    => (others => '0'),
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wvalid    => '0',
    bready    => '0',
    araddr    => (others => '0'),
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arvalid   => '0',
    rready    => '0'
    );

  type at_axil64x40_cmd is array (natural range <>) of rt_axil64x40_cmd;

  --************************************************************************
  --
  --    AXI Lite respone for 64-bit data path and 40-bit addresses.
  --
  --************************************************************************
  type rt_axil64x40_rsp is
  record
    -- Write Address Channel Signals
    awready   : std_logic;
    -- Write Data Channel Signals
    wready    : std_logic;
    -- Write Response Channel
    bresp     : std_logic_vector( 1 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rdata     : std_logic_vector(63 downto 0);
    rresp     : std_logic_vector( 1 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL64x40_RSP_RST     : rt_axil64x40_rsp := (
    awready   => '0',
    wready    => '0',
    bresp     => E_RESP_OKAY,
    bvalid    => '0',
    arready   => '0',
    rdata     => (others => '0'),
    rresp     => E_RESP_OKAY,
    rvalid    => '0'
    );

  type at_axil64x40_rsp is array (natural range <>) of rt_axil64x40_rsp;

  --************************************************************************
  --
  --    AXI Lite command for 64- bit data path and  64 bit addresses.
  --
  --************************************************************************
  type rt_axil64x64_cmd is
  record
    -- Write Address Channel Signals
    awaddr    : std_logic_vector(63 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(63 downto 0);
    wstrb     : std_logic_vector( 7 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    araddr    : std_logic_vector(63 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIL64x64_CMD_RST     : rt_axil64x64_cmd := (
    awaddr    => (others => '0'),
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wvalid    => '0',
    bready    => '0',
    araddr    => (others => '0'),
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arvalid   => '0',
    rready    => '0'
    );

  type at_axil64x64_cmd is array (natural range <>) of rt_axil64x64_cmd;

  --************************************************************************
  --
  -- Even though there is no address bits in the response packets we can hide that detail from the user to make things clearer. We will use alias so that no conversion is needed between
  -- rt_axil64x64_rsp and rt_axil64x32_rsp
  --
  --************************************************************************
  alias rt_axil64x64_rsp    is rt_axil64x32_rsp;
  alias K_AXIL64x64_RSP_RST is K_AXIL64x32_RSP_RST;
  alias at_axil64x64_rsp    is at_axil64x32_rsp;

  --************************************************************************
  --
  --    This is the record AXI Streaming commands from the Master, to the Slave.
  -- It contains all signals sourced by an AXI Stream master and is specifically
  -- for a 16 bit data bus.
  --    If tkeep is always asserted (as in the reset constant), then every transfer
  -- consists of 64-bits of aligned information. This is called a "continuous aligned
  -- stream" and is probably true for most if not all of our AXI Stream Masters.
  --
  --    NOTE: Literally every signal in the AXI streaming protocol is optional. We
  -- implement a subset in these records.
  --
  --************************************************************************
  type rt_axis16_cmd is
  record
    tdata     : std_logic_vector(15 downto 0);  -- primary payload to be transferred to the slave
    tkeep     : std_logic_vector( 1 downto 0);  -- if high the corresponding byte of tdata is to be processed by slave
    tvalid    : std_logic;                      -- high indicates the master desires to transfer tdata to the slave
    tlast     : std_logic;                      -- when asserted it indicates to the slave, the boundary of a packet
    tuser     : std_logic_vector(31 downto 0);  -- Optional user defined signal passed along by AXI interconnect
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIS16_CMD_RST    : rt_axis16_cmd := (
    tdata     => (others => '0'),
    tkeep     => (others => '1'),               -- normally tdata is a "continuous aligned stream"
    tvalid    => '0',
    tlast     => '0',
    tuser     => (others => '0')
    );

  type at_axis16_cmd is array (natural range <>) of rt_axis16_cmd;

  --************************************************************************
  --
  --    The response record for an AXI Stream slave, isn't really much of a
  -- record, but for consistency we'll create a record anyway.
  --
  --************************************************************************
  type rt_axis16_rsp is
  record
    tready    : std_logic;                      -- indicates the slave can accept a transfer in the current clock period
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIS16_RSP_RST   : rt_axis16_rsp := (others => '0');

  type at_axis16_rsp is array (natural range <>) of rt_axis16_rsp;

  -- alternative names
  alias rt_axis32_rsp       is rt_axis16_rsp;
  alias rt_axis64_rsp       is rt_axis16_rsp;
  alias rt_axis128_rsp      is rt_axis16_rsp;
  alias rt_axis256_rsp      is rt_axis16_rsp;
  alias rt_axis512_rsp      is rt_axis16_rsp;
  alias rt_axis1024_rsp     is rt_axis16_rsp;
  alias K_AXIS32_RSP_RST    is K_AXIS16_RSP_RST;
  alias K_AXIS64_RSP_RST    is K_AXIS16_RSP_RST;
  alias K_AXIS128_RSP_RST   is K_AXIS16_RSP_RST;
  alias K_AXIS256_RSP_RST   is K_AXIS16_RSP_RST;
  alias K_AXIS512_RSP_RST   is K_AXIS16_RSP_RST;
  alias K_AXIS1024_RSP_RST  is K_AXIS16_RSP_RST;
  alias at_axis32_rsp       is at_axis16_rsp;
  alias at_axis64_rsp       is at_axis16_rsp;
  alias at_axis128_rsp      is at_axis16_rsp;
  alias at_axis256_rsp      is at_axis16_rsp;
  alias at_axis512_rsp      is at_axis16_rsp;
  alias at_axis1024_rsp     is at_axis16_rsp;

  --************************************************************************
  --
  --    Repeat all these record structures for streaming 32 bit data paths.
  --
  --************************************************************************
  type rt_axis32_cmd is
  record
    tdata     : std_logic_vector(31 downto 0);
    tkeep     : std_logic_vector( 3 downto 0);
    tvalid    : std_logic;
    tlast     : std_logic;
    tuser     : std_logic_vector(31 downto 0);
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIS32_CMD_RST  : rt_axis32_cmd := (
    tdata     => (others => '0'),
    tkeep     => (others => '1'),
    tvalid    => '0',
    tlast     => '0',
    tuser     => (others => '0')
    );

  type at_axis32_cmd is array (natural range <>) of rt_axis32_cmd;

  --************************************************************************
  --
  --    Repeat all these record structures for streaming 64 bit data paths.
  --
  --************************************************************************
  type rt_axis64_cmd is
  record
    tdata     : std_logic_vector(63 downto 0);
    tkeep     : std_logic_vector( 7 downto 0);
    tvalid    : std_logic;
    tlast     : std_logic;
    tuser     : std_logic_vector(31 downto 0);
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIS64_CMD_RST  : rt_axis64_cmd := (
    tdata     => (others => '0'),
    tkeep     => (others => '1'),
    tvalid    => '0',
    tlast     => '0',
    tuser     => (others => '0')
    );

  type at_axis64_cmd is array (natural range <>) of rt_axis64_cmd;

  --************************************************************************
  --
  --    Repeat all these record structures for streaming 128 bit data paths.
  --
  --************************************************************************
  type rt_axis128_cmd is
  record
    tdata     : std_logic_vector(127 downto 0);
    tkeep     : std_logic_vector( 15 downto 0);
    tvalid    : std_logic;
    tlast     : std_logic;
    tuser     : std_logic_vector( 31 downto 0);
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIS128_CMD_RST  : rt_axis128_cmd := (
    tdata     => (others => '0'),
    tkeep     => (others => '1'),
    tvalid    => '0',
    tlast     => '0',
    tuser     => (others => '0')
    );

  type at_axis128_cmd is array (natural range <>) of rt_axis128_cmd;

  --************************************************************************
  --
  --    Repeat all these record structures for streaming 256 bit data paths.
  --
  --************************************************************************
  type rt_axis256_cmd is
  record
    tdata     : std_logic_vector(255 downto 0);
    tkeep     : std_logic_vector( 31 downto 0);
    tvalid    : std_logic;
    tlast     : std_logic;
    tuser     : std_logic_vector( 31 downto 0);
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIS256_CMD_RST  : rt_axis256_cmd := (
    tdata     => (others => '0'),
    tkeep     => (others => '1'),
    tvalid    => '0',
    tlast     => '0',
    tuser     => (others => '0')
    );

  type at_axis256_cmd is array (natural range <>) of rt_axis256_cmd;

  --************************************************************************
  --
  --    Repeat all these record structures for streaming 512 bit data paths.
  --
  --************************************************************************
  type rt_axis512_cmd is
  record
    tdata     : std_logic_vector(511 downto 0);
    tkeep     : std_logic_vector( 63 downto 0);
    tvalid    : std_logic;
    tlast     : std_logic;
    tuser     : std_logic_vector( 31 downto 0);
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIS512_CMD_RST  : rt_axis512_cmd := (
    tdata     => (others => '0'),
    tkeep     => (others => '1'),
    tvalid    => '0',
    tlast     => '0',
    tuser     => (others => '0')
    );

  type at_axis512_cmd is array (natural range <>) of rt_axis512_cmd;

  --************************************************************************
  --
  --    Repeat all these record structures for streaming 1024 bit data paths.
  --
  --************************************************************************
  type rt_axis1024_cmd is
  record
    tdata     : std_logic_vector(1023 downto 0);
    tkeep     : std_logic_vector( 127 downto 0);
    tvalid    : std_logic;
    tlast     : std_logic;
    tuser     : std_logic_vector(  31 downto 0);
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXIS1024_CMD_RST  : rt_axis1024_cmd := (
    tdata     => (others => '0'),
    tkeep     => (others => '1'),
    tvalid    => '0',
    tlast     => '0',
    tuser     => (others => '0')
    );

  type at_axis1024_cmd is array (natural range <>) of rt_axis1024_cmd;


  --************************************************************************
  --
  --    This is the record AXI4 commands from the Master, to the Slave. It
  -- contains all signals sourced by an AXI4 master and is specifically for a
  -- 32 bit data bus and 32 bit address but. These signals are grouped into 5
  -- unique channels as specified by the AXI4 protocol.
  --
  --************************************************************************
  type rt_axi32x32_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector( 7 downto 0);    -- Write addr "tag", all transactions with the same ID bits are responded to in order.
    awaddr    : std_logic_vector(31 downto 0);    -- Write address gives the address of the single transfer
    awlen     : std_logic_vector( 7 downto 0);    -- Burst length gives exact number of transfers in a burst, burst Length = awlen + 1
    awsize    : std_logic_vector( 2 downto 0);    -- Burst size of each transfer in a burst. Bytes=2^awsize (for 64 bits, set awsize="011")
    awburst   : std_logic_vector( 1 downto 0);    -- Burst type and awsize determine how addr for each transfer within the burst is calculated
    awlock    : std_logic_vector( 0 downto 0);    -- Lock type provides additional info about the atomic characteristics of the transfer
    awcache   : std_logic_vector( 3 downto 0);    -- Memory type indicates how transactions progress through a system
    awprot    : std_logic_vector( 2 downto 0);    -- Protection type indicates the privilege and security level
    awqos     : std_logic_vector( 3 downto 0);    -- Quality of Service for each write, "transaction priority" is recommended by the AXI4 spec
    awregion  : std_logic_vector( 3 downto 0);    -- Region id permits a single interface on slave to be used for multiple logical interfaces
    awuser    : std_logic_vector(31 downto 0);    -- Optional user defined signal in the write address channel
    awvalid   : std_logic;                        -- Write address valid, the channel is signaling address and control information
    -- Write Data Channel Signals
    wdata     : std_logic_vector(31 downto 0);    -- Write data
    wstrb     : std_logic_vector( 3 downto 0);    -- Write strobes indicate which byte lanes (in wdata) hold valid data
    wlast     : std_logic;                        -- Write last, this signal indicates the last transfer in a write burst
    wuser     : std_logic_vector(31 downto 0);    -- Optional user defined signal in the write data channel (AXI recommends masters and slaves not use these, but interconnect should support them along A8.3.2)
    wvalid    : std_logic;                        -- Write valid indicates that write data and strobes are available
    -- Write Response Channel
    bready    : std_logic;                        -- Response ready indicates that the master can accept a write response
    -- Read Address Channel
    arid      : std_logic_vector( 7 downto 0);    -- Read addr "tag", AXI4 recommends 4 LSBs for end Masters & 4 MSBs for interconnect Masters
    araddr    : std_logic_vector(31 downto 0);    -- Read address gives the address of the single transfer
    arlen     : std_logic_vector( 7 downto 0);    -- Burst length gives the exact number of transfers in a burst, burst Length = awlen + 1
    arsize    : std_logic_vector( 2 downto 0);    -- Burst size of each transfer in a burst. Bytes=2^arsize (for 64 bits, set arsize = "011")
    arburst   : std_logic_vector( 1 downto 0);    -- Burst type and arsize determine how addr for each transfer within the burst is calculated
    arlock    : std_logic_vector( 0 downto 0);    -- Lock type provides additional info about the atomic characteristics of the transfer
    arcache   : std_logic_vector( 3 downto 0);    -- Memory type indicates how transactions progress through a system
    arprot    : std_logic_vector( 2 downto 0);    -- Protection type, privilege and security level of the transaction
    arqos     : std_logic_vector( 3 downto 0);    -- Quality of Service for each read, "transaction priority" is recommended by the AXI4 spec
    arregion  : std_logic_vector( 3 downto 0);    -- Region id permits a single interface on slave to be used for multiple logical interfaces
    aruser    : std_logic_vector(31 downto 0);    -- Optional user defined signal in the read address channel (AXI recommends masters and slaves not use these, but interconnect should support them along A8.3.2)
    arvalid   : std_logic;                        -- Read address valid, the channel is signaling address and control information
    -- Read Data Channel
    rready    : std_logic;                        -- Read ready indicates the master can accept a read response
  end record;

  -- constant for unconnected or partially connected busses
  constant k_axi32x32_cmd_rst   : rt_axi32x32_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_004BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_004BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi32x32_cmd is array (natural range <>) of rt_axi32x32_cmd;

  --************************************************************************
  --
  --    The record is generated by the slave in response to a previous command.
  -- The direction is "Master In Slave Out", and contains all signals sourced by
  -- an AXI4 slave. These signals are grouped into 5 unique channels as specified
  -- by the AXI4 protocol
  --
  --************************************************************************
  type rt_axi32x32_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;                      -- Write address ready, the slave is ready to accept an address and control signals
    -- Write Data Channel
    wready    : std_logic;                      -- Write ready indicates that the slave can accept the write data
    -- Write Response Channel
    bid       : std_logic_vector( 7 downto 0);  -- Write response ID tag, this signal is the ID tag of the write response
    bresp     : std_logic_vector( 1 downto 0);  -- Write response, indicates the status of the write transaction
    buser     : std_logic_vector(31 downto 0);  -- Optional user defined signal in the write response channel
    bvalid    : std_logic;                      -- Write response valid indicates that the channel is signaling a valid write response
    -- Read Address Channel
    arready   : std_logic;                      -- Read address ready, the slave is ready to accept an address and control signals
    -- Read Data Channel
    rid       : std_logic_vector( 7 downto 0);  -- Read ID tag for the read data group of signals generated by the slave
    rdata     : std_logic_vector(31 downto 0);  -- Read data
    rresp     : std_logic_vector( 1 downto 0);  -- Read response indicates the status of the read transfer
    rlast     : std_logic;                      -- Read last indicates the last transfer in a read burst
    ruser     : std_logic_vector(31 downto 0);  -- Options user defined signal in the read data channel
    rvalid    : std_logic;                      -- Read valid indicates the channel is signaling the requested read data
  end record;

  -- constant for unconnected or partially connected busses
  constant k_axi32x32_rsp_rst    : rt_axi32x32_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi32x32_rsp is array (natural range <>) of rt_axi32x32_rsp;

  --************************************************************************
  --
  --    Repeat all these record structures for 64 bit data paths and 32 bit addresses.
  --
  --************************************************************************
  type rt_axi64x32_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector( 7 downto 0);
    awaddr    : std_logic_vector(31 downto 0);
    awlen     : std_logic_vector( 7 downto 0);
    awsize    : std_logic_vector( 2 downto 0);
    awburst   : std_logic_vector( 1 downto 0);
    awlock    : std_logic_vector( 0 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awqos     : std_logic_vector( 3 downto 0);
    awregion  : std_logic_vector( 3 downto 0);
    awuser    : std_logic_vector(31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(63 downto 0);
    wstrb     : std_logic_vector( 7 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector(31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector( 7 downto 0);
    araddr    : std_logic_vector(31 downto 0);
    arlen     : std_logic_vector( 7 downto 0);
    arsize    : std_logic_vector( 2 downto 0);
    arburst   : std_logic_vector( 1 downto 0);
    arlock    : std_logic_vector( 0 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arqos     : std_logic_vector( 3 downto 0);
    arregion  : std_logic_vector( 3 downto 0);
    aruser    : std_logic_vector(31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI64x32_CMD_RST    : rt_axi64x32_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_008BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_008BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi64x32_cmd is array (natural range <>) of rt_axi64x32_cmd;

  --************************************************************************
  --
  --    Here are 64 bit data, 32 bit address slave responses. (Technically there are no addresses in the response)
  --
  --************************************************************************
  type rt_axi64x32_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector( 7 downto 0);
    bresp     : std_logic_vector( 1 downto 0);
    buser     : std_logic_vector(31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector( 7 downto 0);
    rdata     : std_logic_vector(63 downto 0);
    rresp     : std_logic_vector( 1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector(31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI64x32_RSP_RST    : rt_axi64x32_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi64x32_rsp is array (natural range <>) of rt_axi64x32_rsp;


  --************************************************************************
  --
  --    Repeat all these record structures for 64 bit data paths and 32 bit addresses.
  --
  --************************************************************************
  type rt_axi64x32x16_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector(15 downto 0);
    awaddr    : std_logic_vector(31 downto 0);
    awlen     : std_logic_vector( 7 downto 0);
    awsize    : std_logic_vector( 2 downto 0);
    awburst   : std_logic_vector( 1 downto 0);
    awlock    : std_logic_vector( 0 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awqos     : std_logic_vector( 3 downto 0);
    awregion  : std_logic_vector( 3 downto 0);
    awuser    : std_logic_vector(31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(63 downto 0);
    wstrb     : std_logic_vector( 7 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector(31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector(15 downto 0);
    araddr    : std_logic_vector(31 downto 0);
    arlen     : std_logic_vector( 7 downto 0);
    arsize    : std_logic_vector( 2 downto 0);
    arburst   : std_logic_vector( 1 downto 0);
    arlock    : std_logic_vector( 0 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arqos     : std_logic_vector( 3 downto 0);
    arregion  : std_logic_vector( 3 downto 0);
    aruser    : std_logic_vector(31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI64x32x16_CMD_RST    : rt_axi64x32x16_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_008BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_008BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi64x32x16cmd is array (natural range <>) of rt_axi64x32x16_cmd;

  --************************************************************************
  --
  --    Here are 64 bit data, 32 bit address slave responses. (Technically there are no addresses in the response)
  --
  --************************************************************************
  type rt_axi64x32x16_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector(15 downto 0);
    bresp     : std_logic_vector( 1 downto 0);
    buser     : std_logic_vector(31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector(15 downto 0);
    rdata     : std_logic_vector(63 downto 0);
    rresp     : std_logic_vector( 1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector(31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI64x32x16_RSP_RST    : rt_axi64x32x16_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi64x32x16_rsp is array (natural range <>) of rt_axi64x32x16_rsp;

  --************************************************************************
  --
  --    Here is the command record structures for 512 bit data paths and 32 bit address.
  --
  --************************************************************************
  type rt_axi512x32_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector( 15 downto 0);
    awaddr    : std_logic_vector( 31 downto 0);
    awlen     : std_logic_vector(  7 downto 0);
    awsize    : std_logic_vector(  2 downto 0);
    awburst   : std_logic_vector(  1 downto 0);
    awlock    : std_logic_vector(  0 downto 0);
    awcache   : std_logic_vector(  3 downto 0);
    awprot    : std_logic_vector(  2 downto 0);
    awqos     : std_logic_vector(  3 downto 0);
    awregion  : std_logic_vector(  3 downto 0);
    awuser    : std_logic_vector( 31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(511 downto 0);
    wstrb     : std_logic_vector( 63 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector( 31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector( 15 downto 0);
    araddr    : std_logic_vector( 31 downto 0);
    arlen     : std_logic_vector(  7 downto 0);
    arsize    : std_logic_vector(  2 downto 0);
    arburst   : std_logic_vector(  1 downto 0);
    arlock    : std_logic_vector(  0 downto 0);
    arcache   : std_logic_vector(  3 downto 0);
    arprot    : std_logic_vector(  2 downto 0);
    arqos     : std_logic_vector(  3 downto 0);
    arregion  : std_logic_vector(  3 downto 0);
    aruser    : std_logic_vector( 31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI512X32_CMD_RST   : rt_axi512x32_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_064BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_064BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi512x32_cmd is array (natural range <>) of rt_axi512x32_cmd;

  --************************************************************************
  --
  --    Here are 512 bit slave responses.
  --
  --************************************************************************
  type rt_axi512x32_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector( 15 downto 0);
    bresp     : std_logic_vector(  1 downto 0);
    buser     : std_logic_vector( 31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector( 15 downto 0);
    rdata     : std_logic_vector(511 downto 0);
    rresp     : std_logic_vector(  1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector( 31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI512X32_RSP_RST   : rt_axi512x32_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi512x32_rsp is array (natural range <>) of rt_axi512x32_rsp;


  --************************************************************************
  --
  --    Repeat all these record structures for 128 bit data paths and 40 bit addresses.
  --
  --************************************************************************
  type rt_axi_mpsoc128_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector(15 downto 0);
    awaddr    : std_logic_vector(39 downto 0);
    awlen     : std_logic_vector( 7 downto 0);
    awsize    : std_logic_vector( 2 downto 0);
    awburst   : std_logic_vector( 1 downto 0);
    awlock    : std_logic_vector( 0 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awqos     : std_logic_vector( 3 downto 0);
    awregion  : std_logic_vector( 3 downto 0);
    awuser    : std_logic_vector(15 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(127 downto 0);
    wstrb     : std_logic_vector(15 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector(31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector(15 downto 0);
    araddr    : std_logic_vector(39 downto 0);
    arlen     : std_logic_vector( 7 downto 0);
    arsize    : std_logic_vector( 2 downto 0);
    arburst   : std_logic_vector( 1 downto 0);
    arlock    : std_logic_vector( 0 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arqos     : std_logic_vector( 3 downto 0);
    arregion  : std_logic_vector( 3 downto 0);
    aruser    : std_logic_vector(15 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI_MPSOC128_CMD_RST    : rt_axi_mpsoc128_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_008BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_008BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi_mpsoc128_cmd is array (natural range <>) of rt_axi_mpsoc128_cmd;

  --************************************************************************
  --
  --    Here are 128 bit data, MPSOC 40 bit address slave responses. (Technically there are no addresses in the response)
  --
  --************************************************************************
  type rt_axi_mpsoc128_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector(15 downto 0);
    bresp     : std_logic_vector( 1 downto 0);
    buser     : std_logic_vector(31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector(15 downto 0);
    rdata     : std_logic_vector(127 downto 0);
    rresp     : std_logic_vector( 1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector(31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI_MPSOC128_RSP_RST    : rt_axi_mpsoc128_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi_mpsoc128_rsp is array (natural range <>) of rt_axi_mpsoc128_rsp;


  --************************************************************************
  --
  --    Repeat all these record structures for 64 bit data paths and 40 bit addresses.
  --
  --************************************************************************
  type rt_axi_mpsoc64_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector(15 downto 0);
    awaddr    : std_logic_vector(39 downto 0);
    awlen     : std_logic_vector( 7 downto 0);
    awsize    : std_logic_vector( 2 downto 0);
    awburst   : std_logic_vector( 1 downto 0);
    awlock    : std_logic_vector( 0 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awqos     : std_logic_vector( 3 downto 0);
    awregion  : std_logic_vector( 3 downto 0);
    awuser    : std_logic_vector(15 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(63 downto 0);
    wstrb     : std_logic_vector( 7 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector(31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector(15 downto 0);
    araddr    : std_logic_vector(39 downto 0);
    arlen     : std_logic_vector( 7 downto 0);
    arsize    : std_logic_vector( 2 downto 0);
    arburst   : std_logic_vector( 1 downto 0);
    arlock    : std_logic_vector( 0 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arqos     : std_logic_vector( 3 downto 0);
    arregion  : std_logic_vector( 3 downto 0);
    aruser    : std_logic_vector(15 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI_MPSOC64_CMD_RST    : rt_axi_mpsoc64_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_008BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_008BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi_mpsoc64_cmd is array (natural range <>) of rt_axi_mpsoc64_cmd;

  --************************************************************************
  --
  --    Here are 64 bit data, MPSOC 40 bit address slave responses. (Technically there are no addresses in the response)
  --
  --************************************************************************
  type rt_axi_mpsoc64_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector(15 downto 0);
    bresp     : std_logic_vector( 1 downto 0);
    buser     : std_logic_vector(31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector(15 downto 0);
    rdata     : std_logic_vector(63 downto 0);
    rresp     : std_logic_vector( 1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector(31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI_MPSOC64_RSP_RST    : rt_axi_mpsoc64_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi_mpsoc64_rsp is array (natural range <>) of rt_axi_mpsoc64_rsp;


  --************************************************************************
  --
  --    Repeat all these record structures for 32 bit data paths and MPSOC 40 bit addresses.
  --
  --************************************************************************
  type rt_axi_mpsoc32_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector(15 downto 0);
    awaddr    : std_logic_vector(39 downto 0);
    awlen     : std_logic_vector( 7 downto 0);
    awsize    : std_logic_vector( 2 downto 0);
    awburst   : std_logic_vector( 1 downto 0);
    awlock    : std_logic_vector( 0 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awqos     : std_logic_vector( 3 downto 0);
    awregion  : std_logic_vector( 3 downto 0);
    awuser    : std_logic_vector(15 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(31 downto 0);
    wstrb     : std_logic_vector( 3 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector(31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector(15 downto 0);
    araddr    : std_logic_vector(39 downto 0);
    arlen     : std_logic_vector( 7 downto 0);
    arsize    : std_logic_vector( 2 downto 0);
    arburst   : std_logic_vector( 1 downto 0);
    arlock    : std_logic_vector( 0 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arqos     : std_logic_vector( 3 downto 0);
    arregion  : std_logic_vector( 3 downto 0);
    aruser    : std_logic_vector(15 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI_MPSOC32_CMD_RST    : rt_axi_mpsoc32_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_004BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_004BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi_mpsoc32_cmd is array (natural range <>) of rt_axi_mpsoc32_cmd;

  --************************************************************************
  --
  --    Here are 32 bit data, MPSOC 40 bit address slave responses. (Technically there are no addresses in the response)
  --
  --************************************************************************
  type rt_axi_mpsoc32_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector(15 downto 0);
    bresp     : std_logic_vector( 1 downto 0);
    buser     : std_logic_vector(31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector(15 downto 0);
    rdata     : std_logic_vector(31 downto 0);
    rresp     : std_logic_vector( 1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector(31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI_MPSOC32_RSP_RST    : rt_axi_mpsoc32_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi_mpsoc32_rsp is array (natural range <>) of rt_axi_mpsoc32_rsp;

  --************************************************************************
  --
  --    Repeat all these record structures for 32 bit data paths and 64 bit addresses.
  --
  --************************************************************************
  type rt_axi32_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector( 7 downto 0);
    awaddr    : std_logic_vector(63 downto 0);
    awlen     : std_logic_vector( 7 downto 0);
    awsize    : std_logic_vector( 2 downto 0);
    awburst   : std_logic_vector( 1 downto 0);
    awlock    : std_logic_vector( 0 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awqos     : std_logic_vector( 3 downto 0);
    awregion  : std_logic_vector( 3 downto 0);
    awuser    : std_logic_vector(31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(31 downto 0);
    wstrb     : std_logic_vector( 3 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector(31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector( 7 downto 0);
    araddr    : std_logic_vector(63 downto 0);
    arlen     : std_logic_vector( 7 downto 0);
    arsize    : std_logic_vector( 2 downto 0);
    arburst   : std_logic_vector( 1 downto 0);
    arlock    : std_logic_vector( 0 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arqos     : std_logic_vector( 3 downto 0);
    arregion  : std_logic_vector( 3 downto 0);
    aruser    : std_logic_vector(31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

    -- constant for unconnected or partially connected busses
  constant K_AXI32_CMD_RST    : rt_axi32_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_004BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_004BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi32_cmd is array (natural range <>) of rt_axi32_cmd;

  --************************************************************************
  --
  --    Here are 32 bit data, 64 bit address slave responses. There are no
  -- addresses in the response so we just create an alias to the 32x32 response
  --
  --************************************************************************
  alias rt_axi32_rsp        is rt_axi32x32_rsp;
  alias K_AXI32_RSP_RST     is K_AXI32x32_RSP_RST;
  alias at_axi32_rsp        is at_axi32x32_rsp;

  --************************************************************************
  --
  --    Repeat all these record structures for 64 bit data paths and 64 bit addresses.
  --
  --************************************************************************
  type rt_axi64_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector( 7 downto 0);
    awaddr    : std_logic_vector(63 downto 0);
    awlen     : std_logic_vector( 7 downto 0);
    awsize    : std_logic_vector( 2 downto 0);
    awburst   : std_logic_vector( 1 downto 0);
    awlock    : std_logic_vector( 0 downto 0);
    awcache   : std_logic_vector( 3 downto 0);
    awprot    : std_logic_vector( 2 downto 0);
    awqos     : std_logic_vector( 3 downto 0);
    awregion  : std_logic_vector( 3 downto 0);
    awuser    : std_logic_vector(31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(63 downto 0);
    wstrb     : std_logic_vector( 7 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector(31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector( 7 downto 0);
    araddr    : std_logic_vector(63 downto 0);
    arlen     : std_logic_vector( 7 downto 0);
    arsize    : std_logic_vector( 2 downto 0);
    arburst   : std_logic_vector( 1 downto 0);
    arlock    : std_logic_vector( 0 downto 0);
    arcache   : std_logic_vector( 3 downto 0);
    arprot    : std_logic_vector( 2 downto 0);
    arqos     : std_logic_vector( 3 downto 0);
    arregion  : std_logic_vector( 3 downto 0);
    aruser    : std_logic_vector(31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

    -- constant for unconnected or partially connected busses
  constant K_AXI64_CMD_RST    : rt_axi64_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_008BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_008BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi64_cmd is array (natural range <>) of rt_axi64_cmd;

  --************************************************************************
  --
  --    Here are 64 bit data, 64 bit address slave responses. There are no
  -- addresses in the response so we just create an alias to the 64x32 response
  --
  --************************************************************************
  alias rt_axi64_rsp        is rt_axi64x32_rsp;
  alias K_AXI64_RSP_RST     is K_AXI64x32_RSP_RST;
  alias at_axi64_rsp        is at_axi64x32_rsp;

  --************************************************************************
  --
  --    Repeat all these record structures for 128 bit data paths.
  --
  --************************************************************************
  type rt_axi128_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector(  7 downto 0);
    awaddr    : std_logic_vector( 63 downto 0);
    awlen     : std_logic_vector(  7 downto 0);
    awsize    : std_logic_vector(  2 downto 0);
    awburst   : std_logic_vector(  1 downto 0);
    awlock    : std_logic_vector(  0 downto 0);
    awcache   : std_logic_vector(  3 downto 0);
    awprot    : std_logic_vector(  2 downto 0);
    awqos     : std_logic_vector(  3 downto 0);
    awregion  : std_logic_vector(  3 downto 0);
    awuser    : std_logic_vector( 31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(127 downto 0);
    wstrb     : std_logic_vector( 15 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector( 31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector(  7 downto 0);
    araddr    : std_logic_vector( 63 downto 0);
    arlen     : std_logic_vector(  7 downto 0);
    arsize    : std_logic_vector(  2 downto 0);
    arburst   : std_logic_vector(  1 downto 0);
    arlock    : std_logic_vector(  0 downto 0);
    arcache   : std_logic_vector(  3 downto 0);
    arprot    : std_logic_vector(  2 downto 0);
    arqos     : std_logic_vector(  3 downto 0);
    arregion  : std_logic_vector(  3 downto 0);
    aruser    : std_logic_vector( 31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI128_CMD_RST   : rt_axi128_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_016BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '1',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '1',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_016BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '1'
    );

  type at_axi128_cmd is array (natural range <>) of rt_axi128_cmd;

  --************************************************************************
  --
  --    Here are 128 bit slave responses.
  --
  --************************************************************************
  type rt_axi128_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector(  7 downto 0);
    bresp     : std_logic_vector(  1 downto 0);
    buser     : std_logic_vector( 31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector(  7 downto 0);
    rdata     : std_logic_vector(127 downto 0);
    rresp     : std_logic_vector(  1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector( 31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI128_RSP_RST   : rt_axi128_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi128_rsp is array (natural range <>) of rt_axi128_rsp;

  --************************************************************************
  --
  --    Repeat all these record structures for 256 bit data paths.
  --
  --************************************************************************
  type rt_axi256_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector(  7 downto 0);
    awaddr    : std_logic_vector( 63 downto 0);
    awlen     : std_logic_vector(  7 downto 0);
    awsize    : std_logic_vector(  2 downto 0);
    awburst   : std_logic_vector(  1 downto 0);
    awlock    : std_logic_vector(  0 downto 0);
    awcache   : std_logic_vector(  3 downto 0);
    awprot    : std_logic_vector(  2 downto 0);
    awqos     : std_logic_vector(  3 downto 0);
    awregion  : std_logic_vector(  3 downto 0);
    awuser    : std_logic_vector( 31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(255 downto 0);
    wstrb     : std_logic_vector( 31 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector( 31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector(  7 downto 0);
    araddr    : std_logic_vector( 63 downto 0);
    arlen     : std_logic_vector(  7 downto 0);
    arsize    : std_logic_vector(  2 downto 0);
    arburst   : std_logic_vector(  1 downto 0);
    arlock    : std_logic_vector(  0 downto 0);
    arcache   : std_logic_vector(  3 downto 0);
    arprot    : std_logic_vector(  2 downto 0);
    arqos     : std_logic_vector(  3 downto 0);
    arregion  : std_logic_vector(  3 downto 0);
    aruser    : std_logic_vector( 31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI256_CMD_RST   : rt_axi256_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_032BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_032BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi256_cmd is array (natural range <>) of rt_axi256_cmd;

  --************************************************************************
  --
  --    Here are 256 bit slave responses.
  --
  --************************************************************************
  type rt_axi256_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector(  7 downto 0);
    bresp     : std_logic_vector(  1 downto 0);
    buser     : std_logic_vector( 31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector(  7 downto 0);
    rdata     : std_logic_vector(255 downto 0);
    rresp     : std_logic_vector(  1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector( 31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI256_RSP_RST   : rt_axi256_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '0',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi256_rsp is array (natural range <>) of rt_axi256_rsp;

  --************************************************************************
  --
  --    Here is the command record structures for 512 bit data paths.
  --
  --************************************************************************
  type rt_axi512_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector( 15 downto 0);
    awaddr    : std_logic_vector( 63 downto 0);
    awlen     : std_logic_vector(  7 downto 0);
    awsize    : std_logic_vector(  2 downto 0);
    awburst   : std_logic_vector(  1 downto 0);
    awlock    : std_logic_vector(  0 downto 0);
    awcache   : std_logic_vector(  3 downto 0);
    awprot    : std_logic_vector(  2 downto 0);
    awqos     : std_logic_vector(  3 downto 0);
    awregion  : std_logic_vector(  3 downto 0);
    awuser    : std_logic_vector( 31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(511 downto 0);
    wstrb     : std_logic_vector( 63 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector( 31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector( 15 downto 0);
    araddr    : std_logic_vector( 63 downto 0);
    arlen     : std_logic_vector(  7 downto 0);
    arsize    : std_logic_vector(  2 downto 0);
    arburst   : std_logic_vector(  1 downto 0);
    arlock    : std_logic_vector(  0 downto 0);
    arcache   : std_logic_vector(  3 downto 0);
    arprot    : std_logic_vector(  2 downto 0);
    arqos     : std_logic_vector(  3 downto 0);
    arregion  : std_logic_vector(  3 downto 0);
    aruser    : std_logic_vector( 31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI512_CMD_RST   : rt_axi512_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_064BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '0',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_064BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi512_cmd is array (natural range <>) of rt_axi512_cmd;

    --************************************************************************
  --
  --    Here are 512 bit data, 64 bit address slave responses. There are no
  -- addresses in the response so we just create an alias to the 512x32 response
  --
  --************************************************************************
  alias rt_axi512_rsp        is rt_axi512x32_rsp;
  alias K_AXI512_RSP_RST     is K_AXI512x32_RSP_RST;
  alias at_axi512_rsp        is at_axi512x32_rsp;

  --************************************************************************
  --
  --    Here is the command record structures for 1024 bit data and 64 bit address paths.
  --
  --************************************************************************
  type rt_axi1024_cmd is
  record
    -- Write Address Channel
    awid      : std_logic_vector(   7 downto 0);
    awaddr    : std_logic_vector(  63 downto 0);
    awlen     : std_logic_vector(   7 downto 0);
    awsize    : std_logic_vector(   2 downto 0);
    awburst   : std_logic_vector(   1 downto 0);
    awlock    : std_logic_vector(   0 downto 0);
    awcache   : std_logic_vector(   3 downto 0);
    awprot    : std_logic_vector(   2 downto 0);
    awqos     : std_logic_vector(   3 downto 0);
    awregion  : std_logic_vector(   3 downto 0);
    awuser    : std_logic_vector(  31 downto 0);
    awvalid   : std_logic;
    -- Write Data Channel Signals
    wdata     : std_logic_vector(1023 downto 0);
    wstrb     : std_logic_vector( 127 downto 0);
    wlast     : std_logic;
    wuser     : std_logic_vector(  31 downto 0);
    wvalid    : std_logic;
    -- Write Response Channel
    bready    : std_logic;
    -- Read Address Channel
    arid      : std_logic_vector(   7 downto 0);
    araddr    : std_logic_vector(  63 downto 0);
    arlen     : std_logic_vector(   7 downto 0);
    arsize    : std_logic_vector(   2 downto 0);
    arburst   : std_logic_vector(   1 downto 0);
    arlock    : std_logic_vector(   0 downto 0);
    arcache   : std_logic_vector(   3 downto 0);
    arprot    : std_logic_vector(   2 downto 0);
    arqos     : std_logic_vector(   3 downto 0);
    arregion  : std_logic_vector(   3 downto 0);
    aruser    : std_logic_vector(  31 downto 0);
    arvalid   : std_logic;
    -- Read Data Channel
    rready    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI1024_CMD_RST   : rt_axi1024_cmd := (
    awid      => (others => '0'),
    awaddr    => (others => '0'),
    awlen     => "00000000",
    awsize    => E_SIZE_128BYTES,
    awburst   => E_BURST_INCR,
    awlock    => E_LOCK_NORM,
    awcache   => E_NORM_NCACH_MOD_BUF,
    awprot    => E_NORM_SEC_DATA,
    awqos     => (others => '0'),
    awregion  => (others => '0'),
    awuser    => (others => '0'),
    awvalid   => '0',
    wdata     => (others => '0'),
    wstrb     => (others => '1'),
    wlast     => '1',
    wuser     => (others => '0'),
    wvalid    => '0',
    bready    => '0',
    arid      => (others => '0'),
    araddr    => (others => '0'),
    arlen     => "00000000",
    arsize    => E_SIZE_128BYTES,
    arburst   => E_BURST_INCR,
    arlock    => E_LOCK_NORM,
    arcache   => E_NORM_NCACH_MOD_BUF,
    arprot    => E_NORM_SEC_DATA,
    arqos     => (others => '0'),
    arregion  => (others => '0'),
    aruser    => (others => '0'),
    arvalid   => '0',
    rready    => '0'
    );

  type at_axi1024_cmd is array (natural range <>) of rt_axi1024_cmd;

  --************************************************************************
  --
  --    Here are 1024 bit slave responses.
  --
  --************************************************************************
  type rt_axi1024_rsp is
  record
    -- Write Address Channel
    awready   : std_logic;
    -- Write Data Channel
    wready    : std_logic;
    -- Write Response Channel
    bid       : std_logic_vector(   7 downto 0);
    bresp     : std_logic_vector(   1 downto 0);
    buser     : std_logic_vector(  31 downto 0);
    bvalid    : std_logic;
    -- Read Address Channel
    arready   : std_logic;
    -- Read Data Channel
    rid       : std_logic_vector(   7 downto 0);
    rdata     : std_logic_vector(1023 downto 0);
    rresp     : std_logic_vector(   1 downto 0);
    rlast     : std_logic;
    ruser     : std_logic_vector(  31 downto 0);
    rvalid    : std_logic;
  end record;

  -- constant for unconnected or partially connected busses
  constant K_AXI1024_RSP_RST   : rt_axi1024_rsp := (
    awready  => '0',
    wready   => '0',
    bid      => (others => '0'),
    bresp    => E_RESP_OKAY,
    buser    => (others => '0'),
    bvalid   => '0',
    arready  => '0',
    rid      => (others => '0'),
    rdata    => (others => '0'),
    rresp    => E_RESP_OKAY,
    rlast    => '1',
    ruser    => (others => '0'),
    rvalid   => '0'
    );

  type at_axi1024_rsp is array (natural range <>) of rt_axi1024_rsp;

  --************************************************************************
  --
  --    These are overloaded functions to change AXI command records to/from
  -- 64 bit addressing. When going from 64 to 32 discard MSBs. When going from
  -- 32 to 64, set MSBs to a constant
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axi32x32_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axi32_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axi32_cmd) return  rt_axi32x32_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axi64x32_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axi64_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axi64_cmd) return  rt_axi64x32_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axi512x32_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axi512_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axi512_cmd) return  rt_axi512x32_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axil_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axil32x64_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axil32x64_cmd) return  rt_axil_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axil64x32_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axil64x64_cmd;
  function  axi_addr_resize( i_axi_cmd  : rt_axil64x64_cmd) return  rt_axil64x32_cmd;

end package;

package body axi_pkg is

  --************************************************************************
  --
  -- Upsize the address bits to convert from rt_axi32x32_cmd (32 address bits) to rt_axi32_cmd (64 address bits),
  -- use K_ADDR_MSB as the MSB
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axi32x32_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axi32_cmd is
    variable v_upsized        : rt_axi32_cmd;
  begin
    v_upsized.awid      := i_axi_cmd.awid;
    v_upsized.awaddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.awaddr( 31 downto  0) := i_axi_cmd.awaddr(31 downto 0);
    v_upsized.awlen     := i_axi_cmd.awlen;
    v_upsized.awsize    := i_axi_cmd.awsize;
    v_upsized.awburst   := i_axi_cmd.awburst;
    v_upsized.awlock    := i_axi_cmd.awlock;
    v_upsized.awcache   := i_axi_cmd.awcache;
    v_upsized.awprot    := i_axi_cmd.awprot;
    v_upsized.awqos     := i_axi_cmd.awqos;
    v_upsized.awregion  := i_axi_cmd.awregion;
    v_upsized.awuser    := i_axi_cmd.awuser;
    v_upsized.awvalid   := i_axi_cmd.awvalid;
    v_upsized.wdata     := i_axi_cmd.wdata;
    v_upsized.wstrb     := i_axi_cmd.wstrb;
    v_upsized.wlast     := i_axi_cmd.wlast;
    v_upsized.wuser     := i_axi_cmd.wuser;
    v_upsized.wvalid    := i_axi_cmd.wvalid;
    v_upsized.bready    := i_axi_cmd.bready;
    v_upsized.arid      := i_axi_cmd.arid;
    v_upsized.araddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.araddr( 31 downto  0) := i_axi_cmd.araddr(31 downto 0);
    v_upsized.arlen     := i_axi_cmd.arlen;
    v_upsized.arsize    := i_axi_cmd.arsize;
    v_upsized.arburst   := i_axi_cmd.arburst;
    v_upsized.arlock    := i_axi_cmd.arlock;
    v_upsized.arcache   := i_axi_cmd.arcache;
    v_upsized.arprot    := i_axi_cmd.arprot;
    v_upsized.arqos     := i_axi_cmd.arqos;
    v_upsized.arregion  := i_axi_cmd.arregion;
    v_upsized.aruser    := i_axi_cmd.aruser;
    v_upsized.arvalid   := i_axi_cmd.arvalid;
    v_upsized.rready    := i_axi_cmd.rready;
    return v_upsized;
  end function;

  --************************************************************************
  --
  -- Downsize the address bits to convert from rt_axi32_cmd (64 address bits) to rt_axi32x32_cmd (32 address bits)
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axi32_cmd) return  rt_axi32x32_cmd is
      variable v_downsized      : rt_axi32x32_cmd;
  begin
    v_downsized.awid      := i_axi_cmd.awid;
    v_downsized.awaddr    := i_axi_cmd.awaddr(31 downto 0);
    v_downsized.awlen     := i_axi_cmd.awlen;
    v_downsized.awsize    := i_axi_cmd.awsize;
    v_downsized.awburst   := i_axi_cmd.awburst;
    v_downsized.awlock    := i_axi_cmd.awlock;
    v_downsized.awcache   := i_axi_cmd.awcache;
    v_downsized.awprot    := i_axi_cmd.awprot;
    v_downsized.awqos     := i_axi_cmd.awqos;
    v_downsized.awregion  := i_axi_cmd.awregion;
    v_downsized.awuser    := i_axi_cmd.awuser;
    v_downsized.awvalid   := i_axi_cmd.awvalid;
    v_downsized.wdata     := i_axi_cmd.wdata;
    v_downsized.wstrb     := i_axi_cmd.wstrb;
    v_downsized.wlast     := i_axi_cmd.wlast;
    v_downsized.wuser     := i_axi_cmd.wuser;
    v_downsized.wvalid    := i_axi_cmd.wvalid;
    v_downsized.bready    := i_axi_cmd.bready;
    v_downsized.arid      := i_axi_cmd.arid;
    v_downsized.araddr    := i_axi_cmd.araddr(31 downto 0);
    v_downsized.arlen     := i_axi_cmd.arlen;
    v_downsized.arsize    := i_axi_cmd.arsize;
    v_downsized.arburst   := i_axi_cmd.arburst;
    v_downsized.arlock    := i_axi_cmd.arlock;
    v_downsized.arcache   := i_axi_cmd.arcache;
    v_downsized.arprot    := i_axi_cmd.arprot;
    v_downsized.arqos     := i_axi_cmd.arqos;
    v_downsized.arregion  := i_axi_cmd.arregion;
    v_downsized.aruser    := i_axi_cmd.aruser;
    v_downsized.arvalid   := i_axi_cmd.arvalid;
    v_downsized.rready    := i_axi_cmd.rready;
    return v_downsized;
  end function;

  --************************************************************************
  --
  -- Upsize the address bits to convert from rt_axi64x32_cmd (32 address bits) to rt_axi64_cmd (64 address bits),
  -- use K_ADDR_MSB as the MSB
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axi64x32_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axi64_cmd is
    variable v_upsized        : rt_axi64_cmd;
  begin
    v_upsized.awid      := i_axi_cmd.awid;
    v_upsized.awaddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.awaddr( 31 downto  0) := i_axi_cmd.awaddr(31 downto 0);
    v_upsized.awlen     := i_axi_cmd.awlen;
    v_upsized.awsize    := i_axi_cmd.awsize;
    v_upsized.awburst   := i_axi_cmd.awburst;
    v_upsized.awlock    := i_axi_cmd.awlock;
    v_upsized.awcache   := i_axi_cmd.awcache;
    v_upsized.awprot    := i_axi_cmd.awprot;
    v_upsized.awqos     := i_axi_cmd.awqos;
    v_upsized.awregion  := i_axi_cmd.awregion;
    v_upsized.awuser    := i_axi_cmd.awuser;
    v_upsized.awvalid   := i_axi_cmd.awvalid;
    v_upsized.wdata     := i_axi_cmd.wdata;
    v_upsized.wstrb     := i_axi_cmd.wstrb;
    v_upsized.wlast     := i_axi_cmd.wlast;
    v_upsized.wuser     := i_axi_cmd.wuser;
    v_upsized.wvalid    := i_axi_cmd.wvalid;
    v_upsized.bready    := i_axi_cmd.bready;
    v_upsized.arid      := i_axi_cmd.arid;
    v_upsized.araddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.araddr( 31 downto  0) := i_axi_cmd.araddr(31 downto 0);
    v_upsized.arlen     := i_axi_cmd.arlen;
    v_upsized.arsize    := i_axi_cmd.arsize;
    v_upsized.arburst   := i_axi_cmd.arburst;
    v_upsized.arlock    := i_axi_cmd.arlock;
    v_upsized.arcache   := i_axi_cmd.arcache;
    v_upsized.arprot    := i_axi_cmd.arprot;
    v_upsized.arqos     := i_axi_cmd.arqos;
    v_upsized.arregion  := i_axi_cmd.arregion;
    v_upsized.aruser    := i_axi_cmd.aruser;
    v_upsized.arvalid   := i_axi_cmd.arvalid;
    v_upsized.rready    := i_axi_cmd.rready;
    return v_upsized;
  end function;

  --************************************************************************
  --
  -- Downsize the address bits to convert from rt_axi64_cmd (64 address bits) to rt_axi64x32_cmd (32 address bits)
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axi64_cmd) return  rt_axi64x32_cmd is
    variable v_downsized      : rt_axi64x32_cmd;
  begin
    v_downsized.awid      := i_axi_cmd.awid;
    v_downsized.awaddr    := i_axi_cmd.awaddr(31 downto 0);
    v_downsized.awlen     := i_axi_cmd.awlen;
    v_downsized.awsize    := i_axi_cmd.awsize;
    v_downsized.awburst   := i_axi_cmd.awburst;
    v_downsized.awlock    := i_axi_cmd.awlock;
    v_downsized.awcache   := i_axi_cmd.awcache;
    v_downsized.awprot    := i_axi_cmd.awprot;
    v_downsized.awqos     := i_axi_cmd.awqos;
    v_downsized.awregion  := i_axi_cmd.awregion;
    v_downsized.awuser    := i_axi_cmd.awuser;
    v_downsized.awvalid   := i_axi_cmd.awvalid;
    v_downsized.wdata     := i_axi_cmd.wdata;
    v_downsized.wstrb     := i_axi_cmd.wstrb;
    v_downsized.wlast     := i_axi_cmd.wlast;
    v_downsized.wuser     := i_axi_cmd.wuser;
    v_downsized.wvalid    := i_axi_cmd.wvalid;
    v_downsized.bready    := i_axi_cmd.bready;
    v_downsized.arid      := i_axi_cmd.arid;
    v_downsized.araddr    := i_axi_cmd.araddr(31 downto 0);
    v_downsized.arlen     := i_axi_cmd.arlen;
    v_downsized.arsize    := i_axi_cmd.arsize;
    v_downsized.arburst   := i_axi_cmd.arburst;
    v_downsized.arlock    := i_axi_cmd.arlock;
    v_downsized.arcache   := i_axi_cmd.arcache;
    v_downsized.arprot    := i_axi_cmd.arprot;
    v_downsized.arqos     := i_axi_cmd.arqos;
    v_downsized.arregion  := i_axi_cmd.arregion;
    v_downsized.aruser    := i_axi_cmd.aruser;
    v_downsized.arvalid   := i_axi_cmd.arvalid;
    v_downsized.rready    := i_axi_cmd.rready;
    return v_downsized;
  end function;

  --************************************************************************
  --
  -- Upsize the address bits to convert from rt_axi512x32_cmd (32 address bits) to rt_axi512_cmd (64 address bits),
  -- use K_ADDR_MSB as the MSB
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axi512x32_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axi512_cmd is
    variable v_upsized        : rt_axi512_cmd;
  begin
    v_upsized.awid      := i_axi_cmd.awid;
    v_upsized.awaddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.awaddr( 31 downto  0) := i_axi_cmd.awaddr(31 downto 0);
    v_upsized.awlen     := i_axi_cmd.awlen;
    v_upsized.awsize    := i_axi_cmd.awsize;
    v_upsized.awburst   := i_axi_cmd.awburst;
    v_upsized.awlock    := i_axi_cmd.awlock;
    v_upsized.awcache   := i_axi_cmd.awcache;
    v_upsized.awprot    := i_axi_cmd.awprot;
    v_upsized.awqos     := i_axi_cmd.awqos;
    v_upsized.awregion  := i_axi_cmd.awregion;
    v_upsized.awuser    := i_axi_cmd.awuser;
    v_upsized.awvalid   := i_axi_cmd.awvalid;
    v_upsized.wdata     := i_axi_cmd.wdata;
    v_upsized.wstrb     := i_axi_cmd.wstrb;
    v_upsized.wlast     := i_axi_cmd.wlast;
    v_upsized.wuser     := i_axi_cmd.wuser;
    v_upsized.wvalid    := i_axi_cmd.wvalid;
    v_upsized.bready    := i_axi_cmd.bready;
    v_upsized.arid      := i_axi_cmd.arid;
    v_upsized.araddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.araddr( 31 downto  0) := i_axi_cmd.araddr(31 downto 0);
    v_upsized.arlen     := i_axi_cmd.arlen;
    v_upsized.arsize    := i_axi_cmd.arsize;
    v_upsized.arburst   := i_axi_cmd.arburst;
    v_upsized.arlock    := i_axi_cmd.arlock;
    v_upsized.arcache   := i_axi_cmd.arcache;
    v_upsized.arprot    := i_axi_cmd.arprot;
    v_upsized.arqos     := i_axi_cmd.arqos;
    v_upsized.arregion  := i_axi_cmd.arregion;
    v_upsized.aruser    := i_axi_cmd.aruser;
    v_upsized.arvalid   := i_axi_cmd.arvalid;
    v_upsized.rready    := i_axi_cmd.rready;
    return v_upsized;
  end function;

  --************************************************************************
  --
  -- Downsize the address bits to convert from rt_axi512_cmd (64 address bits) to rt_axi512x32_cmd (32 address bits)
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axi512_cmd) return  rt_axi512x32_cmd is
    variable v_downsized      : rt_axi512x32_cmd;
  begin
    v_downsized.awid      := i_axi_cmd.awid;
    v_downsized.awaddr    := i_axi_cmd.awaddr(31 downto 0);
    v_downsized.awlen     := i_axi_cmd.awlen;
    v_downsized.awsize    := i_axi_cmd.awsize;
    v_downsized.awburst   := i_axi_cmd.awburst;
    v_downsized.awlock    := i_axi_cmd.awlock;
    v_downsized.awcache   := i_axi_cmd.awcache;
    v_downsized.awprot    := i_axi_cmd.awprot;
    v_downsized.awqos     := i_axi_cmd.awqos;
    v_downsized.awregion  := i_axi_cmd.awregion;
    v_downsized.awuser    := i_axi_cmd.awuser;
    v_downsized.awvalid   := i_axi_cmd.awvalid;
    v_downsized.wdata     := i_axi_cmd.wdata;
    v_downsized.wstrb     := i_axi_cmd.wstrb;
    v_downsized.wlast     := i_axi_cmd.wlast;
    v_downsized.wuser     := i_axi_cmd.wuser;
    v_downsized.wvalid    := i_axi_cmd.wvalid;
    v_downsized.bready    := i_axi_cmd.bready;
    v_downsized.arid      := i_axi_cmd.arid;
    v_downsized.araddr    := i_axi_cmd.araddr(31 downto 0);
    v_downsized.arlen     := i_axi_cmd.arlen;
    v_downsized.arsize    := i_axi_cmd.arsize;
    v_downsized.arburst   := i_axi_cmd.arburst;
    v_downsized.arlock    := i_axi_cmd.arlock;
    v_downsized.arcache   := i_axi_cmd.arcache;
    v_downsized.arprot    := i_axi_cmd.arprot;
    v_downsized.arqos     := i_axi_cmd.arqos;
    v_downsized.arregion  := i_axi_cmd.arregion;
    v_downsized.aruser    := i_axi_cmd.aruser;
    v_downsized.arvalid   := i_axi_cmd.arvalid;
    v_downsized.rready    := i_axi_cmd.rready;
    return v_downsized;
  end function;

  --************************************************************************
  --
  -- Upsize the address bits to convert from rt_axil_cmd (32 address bits) to rt_axil32x64_cmd (64 address bits),
  -- use K_ADDR_MSB as the MSB
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axil_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axil32x64_cmd is
    variable v_upsized        : rt_axil32x64_cmd;
  begin
    v_upsized.awaddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.awaddr( 31 downto  0) := i_axi_cmd.awaddr(31 downto 0);
    v_upsized.awcache     := i_axi_cmd.awcache;
    v_upsized.awprot      := i_axi_cmd.awprot ;
    v_upsized.awvalid     := i_axi_cmd.awvalid;
    v_upsized.wdata       := i_axi_cmd.wdata  ;
    v_upsized.wstrb       := i_axi_cmd.wstrb  ;
    v_upsized.wvalid      := i_axi_cmd.wvalid ;
    v_upsized.bready      := i_axi_cmd.bready ;
    v_upsized.araddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.araddr( 31 downto  0) := i_axi_cmd.araddr(31 downto 0);
    v_upsized.arcache     := i_axi_cmd.arcache;
    v_upsized.arprot      := i_axi_cmd.arprot ;
    v_upsized.arvalid     := i_axi_cmd.arvalid;
    v_upsized.rready      := i_axi_cmd.rready ;
    return v_upsized;
  end function;

  --************************************************************************
  --
  -- Downsize the address bits to convert from rt_axil32x64_cmd (64 address bits) to rt_axil_cmd (32 address bits)
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axil32x64_cmd) return  rt_axil_cmd is
    variable v_downsized  : rt_axil_cmd;
  begin
    v_downsized.awaddr    := i_axi_cmd.awaddr(31 downto 0);
    v_downsized.awcache   := i_axi_cmd.awcache;
    v_downsized.awprot    := i_axi_cmd.awprot ;
    v_downsized.awvalid   := i_axi_cmd.awvalid;
    v_downsized.wdata     := i_axi_cmd.wdata  ;
    v_downsized.wstrb     := i_axi_cmd.wstrb  ;
    v_downsized.wvalid    := i_axi_cmd.wvalid ;
    v_downsized.bready    := i_axi_cmd.bready ;
    v_downsized.araddr    := i_axi_cmd.araddr(31 downto 0);
    v_downsized.arcache   := i_axi_cmd.arcache;
    v_downsized.arprot    := i_axi_cmd.arprot ;
    v_downsized.arvalid   := i_axi_cmd.arvalid;
    v_downsized.rready    := i_axi_cmd.rready ;
    return v_downsized;
  end function;

  --************************************************************************
  --
  -- Upsize the address bits to convert from rt_axil64x32_cmd (32 address bits) to rt_axil64x64_cmd (64 address bits),
  -- use K_ADDR_MSB as the MSB
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axil64x32_cmd; K_ADDR_MSB: std_logic_vector(31 downto 0)) return  rt_axil64x64_cmd is
    variable v_upsized        : rt_axil64x64_cmd;
  begin
    v_upsized.awaddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.awaddr( 31 downto  0) := i_axi_cmd.awaddr(31 downto 0);
    v_upsized.awcache     := i_axi_cmd.awcache;
    v_upsized.awprot      := i_axi_cmd.awprot ;
    v_upsized.awvalid     := i_axi_cmd.awvalid;
    v_upsized.wdata       := i_axi_cmd.wdata  ;
    v_upsized.wstrb       := i_axi_cmd.wstrb  ;
    v_upsized.wvalid      := i_axi_cmd.wvalid ;
    v_upsized.bready      := i_axi_cmd.bready ;
    v_upsized.araddr( 63 downto 32) := K_ADDR_MSB;
    v_upsized.araddr( 31 downto  0) := i_axi_cmd.araddr(31 downto 0);
    v_upsized.arcache     := i_axi_cmd.arcache;
    v_upsized.arprot      := i_axi_cmd.arprot ;
    v_upsized.arvalid     := i_axi_cmd.arvalid;
    v_upsized.rready      := i_axi_cmd.rready ;
    return v_upsized;
  end function;

--************************************************************************
  --
  -- Downsize the address bits to convert from rt_axil64x64_cmd (64 address bits) to rt_axil64x32_cmd (32 address bits)
  --
  --************************************************************************
  function  axi_addr_resize( i_axi_cmd  : rt_axil64x64_cmd) return  rt_axil64x32_cmd is
    variable v_downsized  : rt_axil64x32_cmd;
  begin
    v_downsized.awaddr    := i_axi_cmd.awaddr(31 downto 0);
    v_downsized.awcache   := i_axi_cmd.awcache;
    v_downsized.awprot    := i_axi_cmd.awprot ;
    v_downsized.awvalid   := i_axi_cmd.awvalid;
    v_downsized.wdata     := i_axi_cmd.wdata  ;
    v_downsized.wstrb     := i_axi_cmd.wstrb  ;
    v_downsized.wvalid    := i_axi_cmd.wvalid ;
    v_downsized.bready    := i_axi_cmd.bready ;
    v_downsized.araddr    := i_axi_cmd.araddr(31 downto 0);
    v_downsized.arcache   := i_axi_cmd.arcache;
    v_downsized.arprot    := i_axi_cmd.arprot ;
    v_downsized.arvalid   := i_axi_cmd.arvalid;
    v_downsized.rready    := i_axi_cmd.rready ;
    return v_downsized;
  end function;

end package body;
